module machine_jk(
    input wire x,
    input wire CLK,
    input wire RESET,
    output wire F,
    output wire [2:0] S
);

	//jkff jk0(.x(x), .CLK(CLK), .RESET(RESET), .F(), .S());
	//jkff jk1(.x(x), .CLK(CLK), .RESET(RESET), .F(), .S());
	//jkff jk2(.x(x), .CLK(CLK), .RESET(RESET), .F(), .S());


endmodule